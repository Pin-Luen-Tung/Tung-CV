`define CPU_CYCLE     0.7 // 100Mhz
`define MAX           300000000 // 3000000